    Mac OS X            	   2   �                                           ATTR         �   5                  �     com.apple.lastuseddate#PS       �     com.apple.provenance    �     com.dropbox.attrs    ��9g    �[�.     <J����B

f�qͧ��     g�����