    Mac OS X            	   2   �                                           ATTR         �   4                  �     com.apple.lastuseddate#PS       �     com.apple.provenance    �     com.dropbox.attrs    ��2g    EO%     <J����B

f�qͧ��     g���