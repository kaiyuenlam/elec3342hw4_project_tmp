    Mac OS X            	   2   �      �                                      ATTR       �   �   %                  �     com.apple.provenance    �     com.dropbox.attrs     <J����B

f�qͧ��     g��֚�