    Mac OS X            	   2   �                                           ATTR         �   5                  �     com.apple.lastuseddate#PS       �     com.apple.provenance    �     com.dropbox.attrs    �H=g    O�;     )������

f�qͧ��     u���ķ