    Mac OS X            	   2   �                                           ATTR         �   5                  �     com.apple.lastuseddate#PS       �     com.apple.provenance    �     com.dropbox.attrs    ��2g    d�     <J����B

f�qͧ��     g�����