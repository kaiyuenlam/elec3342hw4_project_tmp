    Mac OS X            	   2   �                                           ATTR         �   5                  �     com.apple.lastuseddate#PS       �     com.apple.provenance    �     com.dropbox.attrs    �/2g    �C�     <J����B

f�qͧ��     g��λ�	